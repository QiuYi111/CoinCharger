library verilog;
use verilog.vl_types.all;
entity BtoD_vlg_vec_tst is
end BtoD_vlg_vec_tst;
