library verilog;
use verilog.vl_types.all;
entity D_Controller_vlg_vec_tst is
end D_Controller_vlg_vec_tst;
