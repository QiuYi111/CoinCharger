library verilog;
use verilog.vl_types.all;
entity Translate_vlg_vec_tst is
end Translate_vlg_vec_tst;
