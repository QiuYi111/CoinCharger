library verilog;
use verilog.vl_types.all;
entity scanner_vlg_check_tst is
    port(
        r1              : in     vl_logic;
        r2              : in     vl_logic;
        r3              : in     vl_logic;
        r4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end scanner_vlg_check_tst;
