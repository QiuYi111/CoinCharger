library verilog;
use verilog.vl_types.all;
entity BtoD_vlg_sample_tst is
    port(
        n_0             : in     vl_logic;
        n_1             : in     vl_logic;
        n_2             : in     vl_logic;
        n_3             : in     vl_logic;
        n_4             : in     vl_logic;
        n_5             : in     vl_logic;
        n_6             : in     vl_logic;
        n_7             : in     vl_logic;
        n_8             : in     vl_logic;
        n_9             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end BtoD_vlg_sample_tst;
