library verilog;
use verilog.vl_types.all;
entity scanner_vlg_vec_tst is
end scanner_vlg_vec_tst;
